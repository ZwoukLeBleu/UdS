
*IDEAL:Amplificateur operationnel avec gain boucle ouverte de 100K
.SUBCKT IDEAL 1 2 3
EGAIN 3 0 1 2 1E5
.ENDS
